module testbenchROM();
reg[11:0] A;
wire[7:0] Y;

ROM RR(A, Y);

initial begin
#1
$display("ROM");
$display("A | Y");
$display("-----------|---------");
$monitor("%b |  %b", A, Y);
end
  initial begin
    A = 12'b000000000000;
  #1 A = 12'b000000000001;
  #1 A = 12'b000000000010;
  #1 A = 12'b000000000011;
  #1 A = 12'b000000000100;
  #1 A = 12'b000000000101;
  #1 A = 12'b000000000110;
  #1 A = 12'b000000000111;
  #1 A = 12'b000000001000;
  #1 A = 12'b000000001001;
  #1 A = 12'b000000001010;
  #1 A = 12'b000000001011;
  #1 A = 12'b000000001100;
  #1 A = 12'b000000001101;
  #1 A = 12'b000000001111;
  #1 A = 12'b000000010000;
  #1 A = 12'b000000010001;
  #1 A = 12'b000000010010;
  #1 A = 12'b000000010011;
  #1 A = 12'b000000010100;
  #1 A = 12'b000000010101;
  #1 A = 12'b000000010110;
  #1 A = 12'b000000010111;
  #1 A = 12'b000000011000;





  end

 initial
   #500 $finish;
 initial begin
     $dumpfile("ROM_tb.vcd");
     $dumpvars(0, testbenchROM);
   end
 endmodule
